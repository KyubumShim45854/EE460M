`timescale 1ns / 1ps

module Fitbit();
// HLSM should output to sevenseg : stepcout -> distance covered -> steps over 32(time) -> High activity time


endmodule
